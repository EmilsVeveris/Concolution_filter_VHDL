-- nios2_system_v0.vhd

-- Generated using ACDS version 18.1 625

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity TOP is
	port (
		clk_clk                                                    : in    std_logic                     := '0';             --                              clk.clk
		led_pio_external_connection_export                         : out   std_logic_vector(7 downto 0);                     --      led_pio_external_connection.export
		mem_if_lpddr2_emif_0_pll_ref_clk_clk                       : in    std_logic                     := '0';             -- mem_if_lpddr2_emif_0_pll_ref_clk.clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_mem_clk               : out   std_logic;                                        -- mem_if_lpddr2_emif_0_pll_sharing.pll_mem_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk             : out   std_logic;                                        --                                 .pll_write_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_locked                : out   std_logic;                                        --                                 .pll_locked
		mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk_pre_phy_clk : out   std_logic;                                        --                                 .pll_write_clk_pre_phy_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_addr_cmd_clk          : out   std_logic;                                        --                                 .pll_addr_cmd_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_avl_clk               : out   std_logic;                                        --                                 .pll_avl_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_config_clk            : out   std_logic;                                        --                                 .pll_config_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_mem_phy_clk           : out   std_logic;                                        --                                 .pll_mem_phy_clk
		mem_if_lpddr2_emif_0_pll_sharing_afi_phy_clk               : out   std_logic;                                        --                                 .afi_phy_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_avl_phy_clk           : out   std_logic;                                        --                                 .pll_avl_phy_clk
		mem_if_lpddr2_emif_0_status_local_init_done                : out   std_logic;                                        --      mem_if_lpddr2_emif_0_status.local_init_done
		mem_if_lpddr2_emif_0_status_local_cal_success				  : out   std_logic;                                        --                                 .local_cal_success
		mem_if_lpddr2_emif_0_status_local_cal_fail                 : out   std_logic;                                        --                                 .local_cal_fail
		memory_mem_ca                                              : out   std_logic_vector(9 downto 0);                     --                           memory.mem_ca
		memory_mem_ck                                              : out   std_logic_vector(0 downto 0);                     --                                 .mem_ck
		memory_mem_ck_n                                            : out   std_logic_vector(0 downto 0);                     --                                 .mem_ck_n
		memory_mem_cke                                             : out   std_logic_vector(0 downto 0);                     --                                 .mem_cke
		memory_mem_cs_n                                            : out   std_logic_vector(0 downto 0);                     --                                 .mem_cs_n
		memory_mem_dm                                              : out   std_logic_vector(3 downto 0);                     --                                 .mem_dm
		memory_mem_dq                                              : inout std_logic_vector(31 downto 0) := (others => '0'); --                                 .mem_dq
		memory_mem_dqs                                             : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                 .mem_dqs
		memory_mem_dqs_n                                           : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                 .mem_dqs_n
		oct_rzqin                                                  : in    std_logic                     := '0';             --                              oct.rzqin
		reset_reset_n                                              : in    std_logic                     := '0';             --                            reset.reset_n                   --    seg_pio_2_external_connection.export
		sw_pio_external_connection_export                          : in    std_logic_vector(7 downto 0)  := (others => '0'); --       sw_pio_external_connection.export
		uart_0_external_connection_rxd                             : in    std_logic                     := '0';             --       uart_0_external_connection.rxd
		uart_0_external_connection_txd                             : out   std_logic;                                        --                                 .txd
				
		I2C_SCL : inout std_logic;
		
		I2C_SDA : inout std_logic;

		HDMI_TX_CLK : out std_logic;
		HDMI_TX_D : out std_logic_vector(23 downto 0);
		HDMI_TX_DE : out std_logic;
		HDMI_TX_HS : out std_logic;
		HDMI_TX_INT : in std_logic;
		HDMI_TX_VS : buffer std_logic

	);
end entity TOP;


architecture behavioral of TOP is

	component nios2_system_v0 is
	port (
		clk_clk                                                    : in    std_logic                     := '0';             --                              clk.clk
		data_out_external_connection_export                        : out   std_logic_vector(7 downto 0);                    --     data_out_external_connection.export
		led_pio_external_connection_export                         : out   std_logic_vector(7 downto 0);                     --      led_pio_external_connection.export
		mem_if_lpddr2_emif_0_pll_sharing_pll_mem_clk               : out   std_logic;                                        -- mem_if_lpddr2_emif_0_pll_sharing.pll_mem_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk             : out   std_logic;                                        --                                 .pll_write_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_locked                : out   std_logic;                                        --                                 .pll_locked
		mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk_pre_phy_clk : out   std_logic;                                        --                                 .pll_write_clk_pre_phy_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_addr_cmd_clk          : out   std_logic;                                        --                                 .pll_addr_cmd_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_avl_clk               : out   std_logic;                                        --                                 .pll_avl_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_config_clk            : out   std_logic;                                        --                                 .pll_config_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_mem_phy_clk           : out   std_logic;                                        --                                 .pll_mem_phy_clk
		mem_if_lpddr2_emif_0_pll_sharing_afi_phy_clk               : out   std_logic;                                        --                                 .afi_phy_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_avl_phy_clk           : out   std_logic;                                        --                                 .pll_avl_phy_clk
		mem_if_lpddr2_emif_0_status_local_init_done                : out   std_logic;                                        --      mem_if_lpddr2_emif_0_status.local_init_done
		mem_if_lpddr2_emif_0_status_local_cal_success              : out   std_logic;                                        --                                 .local_cal_success
		mem_if_lpddr2_emif_0_status_local_cal_fail                 : out   std_logic;                                        --                                 .local_cal_fail
		memory_mem_ca                                              : out   std_logic_vector(9 downto 0);                     --                           memory.mem_ca
		memory_mem_ck                                              : out   std_logic_vector(0 downto 0);                     --                                 .mem_ck
		memory_mem_ck_n                                            : out   std_logic_vector(0 downto 0);                     --                                 .mem_ck_n
		memory_mem_cke                                             : out   std_logic_vector(0 downto 0);                     --                                 .mem_cke
		memory_mem_cs_n                                            : out   std_logic_vector(0 downto 0);                     --                                 .mem_cs_n
		memory_mem_dm                                              : out   std_logic_vector(3 downto 0);                     --                                 .mem_dm
		memory_mem_dq                                              : inout std_logic_vector(31 downto 0) := (others => '0'); --                                 .mem_dq
		memory_mem_dqs                                             : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                 .mem_dqs
		memory_mem_dqs_n                                           : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                 .mem_dqs_n
		oct_rzqin                                                  : in    std_logic                     := '0';             --                              oct.rzqin
		reset_reset_n                                              : in    std_logic                     := '0';             --                            reset.reset_n
		start_bit_external_connection_export                       : out   std_logic;
		sw_pio_external_connection_export                          : in    std_logic_vector(7 downto 0)  := (others => '0'); --       sw_pio_external_connection.export
		uart_0_external_connection_rxd                             : in    std_logic                     := '0';             --       uart_0_external_connection.rxd
		uart_0_external_connection_txd                             : out   std_logic;                                        --                                 .txd
		write_en_external_connection_export                        : out   std_logic;  
		reset_cnt_external_connection_export                       : out   std_logic
	);
	end component;
	
		component periphery_ctrl is
		generic
		(
			CLK_SPEED : integer := 50_000_000
		);
		port
		(
			i_clk : in std_logic;
			i_reset_n : in std_logic := '1';
			i_int_n : in std_logic := '1';
			io_sda : inout std_logic;
			io_scl : inout std_logic;
			o_status : out std_logic_vector(7 downto 0);
			o_ack_error : out std_logic
		);
	end component;
	
		component COUNTER_GEN_1 is
	generic(
				WIDTH: integer  :=	8
	);
	port (
		 RESET_N,CLK,EN,CLC,DIR : IN std_logic;
		 CNT : OUT std_logic_vector(WIDTH-1 downto 0)
	);
	end component;
	

signal s_ack_error : std_logic;
signal HDMI_DEN_net : std_logic;
signal ClkDividerCntOut : std_logic_vector(22 downto 0);
signal cpu_data, ram_data : std_logic_vector(7 downto 0);
signal fsm_en : std_logic;
signal address, RAM_ADDR : std_logic_vector(18 downto 0);
signal Enable : std_logic;
signal R_IN_net,G_IN_net,B_IN_net : std_logic_vector(7 downto 0);

SIGNAL X_cord : std_logic_vector(9 downto 0);
SIGNAL Y_cord : std_logic_vector(9 downto 0);
signal RESET_CNT, wren, REC_DATA, Start_bit : std_logic;
	
begin	
	
	   VGA_DRIVER : entity work.VGA_DRIVER
	generic map
	(
		H_FP => 16,
		H_PULSE => 96,
		H_BP => 48,
		H_PIXELS => 640,
		V_FP => 10,
		V_PULSE => 2,
		V_BP => 29,
		V_PIXELS => 480
	)
	port map
	(
		RESET_N => reset_reset_n,
		CLK => ClkDividerCntOut(0),
		EN => '1',
		X => X_cord,
		Y => y_cord,
		
		R_IN =>R_IN_net,
	   G_IN =>G_IN_net,
	   B_IN =>B_IN_net,
	
		HDMI_TX_D => HDMI_TX_D,
		HDMI_DEN => HDMI_TX_DE,
		HDMI_VSYNC => HDMI_TX_VS,
		HDMI_HSYNC => HDMI_TX_HS
	);
NIOS_2 : nios2_system_v0 port map
(
		clk_clk => clk_clk,
		data_out_external_connection_export										=> cpu_data,
		led_pio_external_connection_export 										=> led_pio_external_connection_export,
		mem_if_lpddr2_emif_0_pll_sharing_pll_mem_clk							=> mem_if_lpddr2_emif_0_pll_sharing_pll_mem_clk,
		mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk                 => mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk,
		mem_if_lpddr2_emif_0_pll_sharing_pll_locked							=> mem_if_lpddr2_emif_0_pll_sharing_pll_locked,
		mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk_pre_phy_clk		=> mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk_pre_phy_clk,
		mem_if_lpddr2_emif_0_pll_sharing_pll_addr_cmd_clk					=> mem_if_lpddr2_emif_0_pll_sharing_pll_addr_cmd_clk,
		mem_if_lpddr2_emif_0_pll_sharing_pll_avl_clk							=> mem_if_lpddr2_emif_0_pll_sharing_pll_avl_clk,
		mem_if_lpddr2_emif_0_pll_sharing_pll_config_clk						=> mem_if_lpddr2_emif_0_pll_sharing_pll_config_clk,
		mem_if_lpddr2_emif_0_pll_sharing_pll_mem_phy_clk					=> mem_if_lpddr2_emif_0_pll_sharing_pll_mem_phy_clk,
		mem_if_lpddr2_emif_0_pll_sharing_afi_phy_clk							=> mem_if_lpddr2_emif_0_pll_sharing_afi_phy_clk,
		mem_if_lpddr2_emif_0_pll_sharing_pll_avl_phy_clk					=> mem_if_lpddr2_emif_0_pll_sharing_pll_avl_phy_clk,
		mem_if_lpddr2_emif_0_status_local_init_done							=> mem_if_lpddr2_emif_0_status_local_init_done,
		mem_if_lpddr2_emif_0_status_local_cal_success						=> mem_if_lpddr2_emif_0_status_local_cal_success,
		mem_if_lpddr2_emif_0_status_local_cal_fail  							=> mem_if_lpddr2_emif_0_status_local_cal_fail, 
		memory_mem_ca																	=> memory_mem_ca,
		memory_mem_ck																	=> memory_mem_ck,
		memory_mem_ck_n																=> memory_mem_ck_n,
		memory_mem_cke																	=> memory_mem_cke,
		memory_mem_cs_n																=> memory_mem_cs_n,
		memory_mem_dm																	=> memory_mem_dm,
		memory_mem_dq																	=> memory_mem_dq,
		memory_mem_dqs																	=> memory_mem_dqs,
		memory_mem_dqs_n 																=> memory_mem_dqs_n,
		oct_rzqin																		=> oct_rzqin,	
		reset_reset_n 																	=> reset_reset_n,
		sw_pio_external_connection_export 										=> sw_pio_external_connection_export,
		uart_0_external_connection_rxd											=> uart_0_external_connection_rxd,
		uart_0_external_connection_txd											=> uart_0_external_connection_txd,
		write_en_external_connection_export										=> REC_DATA,
		start_bit_external_connection_export									=> Start_bit,
		reset_cnt_external_connection_export                       		=> RESET_CNT
		);
		
	pc : periphery_ctrl port map
	(
		i_clk => clk_clk,
		i_reset_n => reset_reset_n,
		i_int_n => HDMI_TX_INT,
		io_sda => I2C_SDA,
		io_scl => I2C_SCL,
		o_status => open,
		o_ack_error => s_ack_error
	);

	CNT_ADDR : entity work.COUNTER_GEN_1
		generic map(WIDTH => 19)
		port map (
			RESET_N => HDMI_TX_VS,
			CLK => ClkDividerCntOut(0),
			EN => Enable,
			CLC=> '0',
			DIR => '1',
			CNT => address
			);
			
	CNT_WRITE_ADDR : entity work.COUNTER_GEN_1
		generic map(WIDTH => 19)
		port map (
			RESET_N => RESET_CNT,
			CLK => clk_clk,
			EN => fsm_en,
			CLC=> '0',
			DIR => '1',
			CNT => RAM_ADDR
			);
			
		CLK_DIVIDER : COUNTER_GEN_1
		generic map(WIDTH => 23)
		port map (RESET_N => reset_reset_n,
					 CLK => clk_clk,
					 EN => reset_reset_n,
					 CLC=> '0',
					 DIR => '1',
					 CNT => ClkDividerCntOut
	);

RAM_0 : entity work.RAM_0
	port map (
		clock => clk_clk,
		data => cpu_data, 
		rdaddress => address,
		wraddress => RAM_ADDR,
		wren =>wren,
		q => ram_data
	);
	FSM_RECIVE : entity work.FSM_RECIVE
		port map (
		CLK => clk_clk,
		RESET_N => reset_reset_n,
		REC_DATA => REC_DATA, 
		WREN => wren,
		CNT_EN => fsm_en,
		Start_bit => Start_bit
	);
	
		Blue_Square: process(X_cord,Y_cord)
	begin
	
		if (X_cord < 640) and (Y_cord < 480) then
						R_IN_net <= ram_data;
						G_IN_net <= ram_data;
						B_IN_net <= ram_data;
						Enable <= '1';

		else
						R_IN_net <= (others => '0');
						G_IN_net <= (others => '1');
						B_IN_net <= (others => '0');
						Enable <= '0';

		end if;
	end process;

	HDMI_TX_CLK <= ClkDividerCntOut(0);
--	HDMI_TX_DE <= HDMI_DEN_net;

	
end;
