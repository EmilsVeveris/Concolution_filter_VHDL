-- nios2_system_v0.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios2_system_v0 is
	port (
		audio_0_external_interface_ADCDAT    : in  std_logic                    := '0';             --    audio_0_external_interface.ADCDAT
		audio_0_external_interface_ADCLRCK   : in  std_logic                    := '0';             --                              .ADCLRCK
		audio_0_external_interface_BCLK      : in  std_logic                    := '0';             --                              .BCLK
		audio_0_external_interface_DACDAT    : out std_logic;                                       --                              .DACDAT
		audio_0_external_interface_DACLRCK   : in  std_logic                    := '0';             --                              .DACLRCK
		audio_xclk_clk                       : out std_logic;                                       --                    audio_xclk.clk
		clk_clk                              : in  std_logic                    := '0';             --                           clk.clk
		i2c_0_i2c_serial_sda_inout           : inout  std_logic                    := '0';             --              i2c_0_i2c_serial.sda_in
		i2c_0_i2c_serial_scl_inout           : inout  std_logic                    := '0';             --                              .scl_in

		led_pio_external_connection_export   : out std_logic_vector(7 downto 0);                    --   led_pio_external_connection.export
		reset_reset_n                        : in  std_logic                    := '0';             --                         reset.reset_n
		seg_pio_0_external_connection_export : out std_logic_vector(7 downto 0);                    -- seg_pio_0_external_connection.export
		seg_pio_1_external_connection_export : out std_logic_vector(7 downto 0);                    -- seg_pio_1_external_connection.export
		seg_pio_2_external_connection_export : out std_logic_vector(7 downto 0);                    -- seg_pio_2_external_connection.export
		sw_pio_external_connection_export    : in  std_logic_vector(7 downto 0) := (others => '0')  --    sw_pio_external_connection.export
	);
end entity nios2_system_v0;

architecture rtl of nios2_system_v0 is
	component nios2_system_v0_audio_0 is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			read        : in  std_logic                     := 'X';             -- read
			write       : in  std_logic                     := 'X';             -- write
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			irq         : out std_logic;                                        -- irq
			AUD_ADCDAT  : in  std_logic                     := 'X';             -- export
			AUD_ADCLRCK : in  std_logic                     := 'X';             -- export
			AUD_BCLK    : in  std_logic                     := 'X';             -- export
			AUD_DACDAT  : out std_logic;                                        -- export
			AUD_DACLRCK : in  std_logic                     := 'X'              -- export
		);
	end component nios2_system_v0_audio_0;

	component nios2_system_v0_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(16 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(16 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component nios2_system_v0_cpu;

	component altera_avalon_i2c is
		generic (
			USE_AV_ST       : integer := 0;
			FIFO_DEPTH      : integer := 4;
			FIFO_DEPTH_LOG2 : integer := 2
		);
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			rst_n     : in  std_logic                     := 'X';             -- reset_n
			intr      : out std_logic;                                        -- irq
			addr      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			sda_in    : in  std_logic                     := 'X';             -- sda_in
			scl_in    : in  std_logic                     := 'X';             -- scl_in
			sda_oe    : out std_logic;                                        -- sda_oe
			scl_oe    : out std_logic;                                        -- scl_oe
			src_data  : out std_logic_vector(7 downto 0);                     -- data
			src_valid : out std_logic;                                        -- valid
			src_ready : in  std_logic                     := 'X';             -- ready
			snk_data  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			snk_valid : in  std_logic                     := 'X';             -- valid
			snk_ready : out std_logic                                         -- ready
		);
	end component altera_avalon_i2c;

	component nios2_system_v0_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios2_system_v0_jtag_uart;

	component nios2_system_v0_led_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component nios2_system_v0_led_pio;

	component nios2_system_v0_onchip_mem is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component nios2_system_v0_onchip_mem;

	component nios2_system_v0_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component nios2_system_v0_pll_0;

	component nios2_system_v0_sw_pio is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component nios2_system_v0_sw_pio;

	component nios2_system_v0_sys_clk_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios2_system_v0_sys_clk_timer;

	component nios2_system_v0_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component nios2_system_v0_sysid;

	component nios2_system_v0_mm_interconnect_0 is
		port (
			clk_0_clk_clk                             : in  std_logic                     := 'X';             -- clk
			pll_0_outclk0_clk                         : in  std_logic                     := 'X';             -- clk
			audio_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			cpu_reset_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                   : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest               : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                      : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                     : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess               : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address            : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest        : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read               : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_instruction_master_readdatavalid      : out std_logic;                                        -- readdatavalid
			audio_0_avalon_audio_slave_address        : out std_logic_vector(1 downto 0);                     -- address
			audio_0_avalon_audio_slave_write          : out std_logic;                                        -- write
			audio_0_avalon_audio_slave_read           : out std_logic;                                        -- read
			audio_0_avalon_audio_slave_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_0_avalon_audio_slave_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			audio_0_avalon_audio_slave_chipselect     : out std_logic;                                        -- chipselect
			cpu_debug_mem_slave_address               : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write                 : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                  : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess           : out std_logic;                                        -- debugaccess
			i2c_0_csr_address                         : out std_logic_vector(3 downto 0);                     -- address
			i2c_0_csr_write                           : out std_logic;                                        -- write
			i2c_0_csr_read                            : out std_logic;                                        -- read
			i2c_0_csr_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i2c_0_csr_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_address       : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write         : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read          : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect    : out std_logic;                                        -- chipselect
			led_pio_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			led_pio_s1_write                          : out std_logic;                                        -- write
			led_pio_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_pio_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			led_pio_s1_chipselect                     : out std_logic;                                        -- chipselect
			onchip_mem_s1_address                     : out std_logic_vector(12 downto 0);                    -- address
			onchip_mem_s1_write                       : out std_logic;                                        -- write
			onchip_mem_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_mem_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_mem_s1_byteenable                  : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_mem_s1_chipselect                  : out std_logic;                                        -- chipselect
			onchip_mem_s1_clken                       : out std_logic;                                        -- clken
			seg_pio_0_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			seg_pio_0_s1_write                        : out std_logic;                                        -- write
			seg_pio_0_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			seg_pio_0_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			seg_pio_0_s1_chipselect                   : out std_logic;                                        -- chipselect
			seg_pio_1_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			seg_pio_1_s1_write                        : out std_logic;                                        -- write
			seg_pio_1_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			seg_pio_1_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			seg_pio_1_s1_chipselect                   : out std_logic;                                        -- chipselect
			seg_pio_2_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			seg_pio_2_s1_write                        : out std_logic;                                        -- write
			seg_pio_2_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			seg_pio_2_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			seg_pio_2_s1_chipselect                   : out std_logic;                                        -- chipselect
			sw_pio_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			sw_pio_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sys_clk_timer_s1_address                  : out std_logic_vector(2 downto 0);                     -- address
			sys_clk_timer_s1_write                    : out std_logic;                                        -- write
			sys_clk_timer_s1_readdata                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sys_clk_timer_s1_writedata                : out std_logic_vector(15 downto 0);                    -- writedata
			sys_clk_timer_s1_chipselect               : out std_logic;                                        -- chipselect
			sysid_control_slave_address               : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component nios2_system_v0_mm_interconnect_0;

	component nios2_system_v0_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios2_system_v0_irq_mapper;

	component nios2_system_v0_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios2_system_v0_rst_controller;

	component nios2_system_v0_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios2_system_v0_rst_controller_001;

	signal pll_0_outclk0_clk                                             : std_logic;                     -- pll_0:outclk_0 -> [audio_xclk_clk, audio_0:clk, mm_interconnect_0:pll_0_outclk0_clk, rst_controller:clk]
	signal cpu_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                   : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                       : std_logic_vector(16 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                          : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_write                                         : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                     : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                : std_logic_vector(16 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                   : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal cpu_instruction_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	signal mm_interconnect_0_audio_0_avalon_audio_slave_chipselect       : std_logic;                     -- mm_interconnect_0:audio_0_avalon_audio_slave_chipselect -> audio_0:chipselect
	signal mm_interconnect_0_audio_0_avalon_audio_slave_readdata         : std_logic_vector(31 downto 0); -- audio_0:readdata -> mm_interconnect_0:audio_0_avalon_audio_slave_readdata
	signal mm_interconnect_0_audio_0_avalon_audio_slave_address          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_0_avalon_audio_slave_address -> audio_0:address
	signal mm_interconnect_0_audio_0_avalon_audio_slave_read             : std_logic;                     -- mm_interconnect_0:audio_0_avalon_audio_slave_read -> audio_0:read
	signal mm_interconnect_0_audio_0_avalon_audio_slave_write            : std_logic;                     -- mm_interconnect_0:audio_0_avalon_audio_slave_write -> audio_0:write
	signal mm_interconnect_0_audio_0_avalon_audio_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_0_avalon_audio_slave_writedata -> audio_0:writedata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                 : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_i2c_0_csr_readdata                          : std_logic_vector(31 downto 0); -- i2c_0:readdata -> mm_interconnect_0:i2c_0_csr_readdata
	signal mm_interconnect_0_i2c_0_csr_address                           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:i2c_0_csr_address -> i2c_0:addr
	signal mm_interconnect_0_i2c_0_csr_read                              : std_logic;                     -- mm_interconnect_0:i2c_0_csr_read -> i2c_0:read
	signal mm_interconnect_0_i2c_0_csr_write                             : std_logic;                     -- mm_interconnect_0:i2c_0_csr_write -> i2c_0:write
	signal mm_interconnect_0_i2c_0_csr_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:i2c_0_csr_writedata -> i2c_0:writedata
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest             : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_mem_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_chipselect -> onchip_mem:chipselect
	signal mm_interconnect_0_onchip_mem_s1_readdata                      : std_logic_vector(31 downto 0); -- onchip_mem:readdata -> mm_interconnect_0:onchip_mem_s1_readdata
	signal mm_interconnect_0_onchip_mem_s1_address                       : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_mem_s1_address -> onchip_mem:address
	signal mm_interconnect_0_onchip_mem_s1_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_mem_s1_byteenable -> onchip_mem:byteenable
	signal mm_interconnect_0_onchip_mem_s1_write                         : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_write -> onchip_mem:write
	signal mm_interconnect_0_onchip_mem_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_mem_s1_writedata -> onchip_mem:writedata
	signal mm_interconnect_0_onchip_mem_s1_clken                         : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_clken -> onchip_mem:clken
	signal mm_interconnect_0_sys_clk_timer_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	signal mm_interconnect_0_sys_clk_timer_s1_readdata                   : std_logic_vector(15 downto 0); -- sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	signal mm_interconnect_0_sys_clk_timer_s1_address                    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	signal mm_interconnect_0_sys_clk_timer_s1_write                      : std_logic;                     -- mm_interconnect_0:sys_clk_timer_s1_write -> mm_interconnect_0_sys_clk_timer_s1_write:in
	signal mm_interconnect_0_sys_clk_timer_s1_writedata                  : std_logic_vector(15 downto 0); -- mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	signal mm_interconnect_0_led_pio_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:led_pio_s1_chipselect -> led_pio:chipselect
	signal mm_interconnect_0_led_pio_s1_readdata                         : std_logic_vector(31 downto 0); -- led_pio:readdata -> mm_interconnect_0:led_pio_s1_readdata
	signal mm_interconnect_0_led_pio_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_pio_s1_address -> led_pio:address
	signal mm_interconnect_0_led_pio_s1_write                            : std_logic;                     -- mm_interconnect_0:led_pio_s1_write -> mm_interconnect_0_led_pio_s1_write:in
	signal mm_interconnect_0_led_pio_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_pio_s1_writedata -> led_pio:writedata
	signal mm_interconnect_0_seg_pio_0_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:seg_pio_0_s1_chipselect -> seg_pio_0:chipselect
	signal mm_interconnect_0_seg_pio_0_s1_readdata                       : std_logic_vector(31 downto 0); -- seg_pio_0:readdata -> mm_interconnect_0:seg_pio_0_s1_readdata
	signal mm_interconnect_0_seg_pio_0_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:seg_pio_0_s1_address -> seg_pio_0:address
	signal mm_interconnect_0_seg_pio_0_s1_write                          : std_logic;                     -- mm_interconnect_0:seg_pio_0_s1_write -> mm_interconnect_0_seg_pio_0_s1_write:in
	signal mm_interconnect_0_seg_pio_0_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:seg_pio_0_s1_writedata -> seg_pio_0:writedata
	signal mm_interconnect_0_seg_pio_1_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:seg_pio_1_s1_chipselect -> seg_pio_1:chipselect
	signal mm_interconnect_0_seg_pio_1_s1_readdata                       : std_logic_vector(31 downto 0); -- seg_pio_1:readdata -> mm_interconnect_0:seg_pio_1_s1_readdata
	signal mm_interconnect_0_seg_pio_1_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:seg_pio_1_s1_address -> seg_pio_1:address
	signal mm_interconnect_0_seg_pio_1_s1_write                          : std_logic;                     -- mm_interconnect_0:seg_pio_1_s1_write -> mm_interconnect_0_seg_pio_1_s1_write:in
	signal mm_interconnect_0_seg_pio_1_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:seg_pio_1_s1_writedata -> seg_pio_1:writedata
	signal mm_interconnect_0_seg_pio_2_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:seg_pio_2_s1_chipselect -> seg_pio_2:chipselect
	signal mm_interconnect_0_seg_pio_2_s1_readdata                       : std_logic_vector(31 downto 0); -- seg_pio_2:readdata -> mm_interconnect_0:seg_pio_2_s1_readdata
	signal mm_interconnect_0_seg_pio_2_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:seg_pio_2_s1_address -> seg_pio_2:address
	signal mm_interconnect_0_seg_pio_2_s1_write                          : std_logic;                     -- mm_interconnect_0:seg_pio_2_s1_write -> mm_interconnect_0_seg_pio_2_s1_write:in
	signal mm_interconnect_0_seg_pio_2_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:seg_pio_2_s1_writedata -> seg_pio_2:writedata
	signal mm_interconnect_0_sw_pio_s1_readdata                          : std_logic_vector(31 downto 0); -- sw_pio:readdata -> mm_interconnect_0:sw_pio_s1_readdata
	signal mm_interconnect_0_sw_pio_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sw_pio_s1_address -> sw_pio:address
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- sys_clk_timer:irq -> irq_mapper:receiver1_irq
	signal cpu_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [audio_0:reset, mm_interconnect_0:audio_0_reset_reset_bridge_in_reset_reset]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_mem:reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_001_reset_out_reset_req                        : std_logic;                     -- rst_controller_001:reset_req -> [cpu:reset_req, onchip_mem:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> [pll_0:rst, rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_sys_clk_timer_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_0_sys_clk_timer_s1_write:inv -> sys_clk_timer:write_n
	signal mm_interconnect_0_led_pio_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_led_pio_s1_write:inv -> led_pio:write_n
	signal mm_interconnect_0_seg_pio_0_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_seg_pio_0_s1_write:inv -> seg_pio_0:write_n
	signal mm_interconnect_0_seg_pio_1_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_seg_pio_1_s1_write:inv -> seg_pio_1:write_n
	signal mm_interconnect_0_seg_pio_2_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_seg_pio_2_s1_write:inv -> seg_pio_2:write_n
	signal rst_controller_001_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [cpu:reset_n, i2c_0:rst_n, jtag_uart:rst_n, led_pio:reset_n, seg_pio_0:reset_n, seg_pio_1:reset_n, seg_pio_2:reset_n, sw_pio:reset_n, sys_clk_timer:reset_n, sysid:reset_n]
	
	signal I2C_DIN_net, I2C_CLK_net : std_logic;
	signal I2C_SERIAL_SDA_IN_net, I2C_SERIAL_SCL_IN_net : std_logic;
	signal I2C_SERIAL_SDA_OE_net, I2C_SERIAL_SCL_OE_net : std_logic;
	
begin

	audio_0 : component nios2_system_v0_audio_0
		port map (
			clk         => pll_0_outclk0_clk,                                       --                clk.clk
			reset       => rst_controller_reset_out_reset,                          --              reset.reset
			address     => mm_interconnect_0_audio_0_avalon_audio_slave_address,    -- avalon_audio_slave.address
			chipselect  => mm_interconnect_0_audio_0_avalon_audio_slave_chipselect, --                   .chipselect
			read        => mm_interconnect_0_audio_0_avalon_audio_slave_read,       --                   .read
			write       => mm_interconnect_0_audio_0_avalon_audio_slave_write,      --                   .write
			writedata   => mm_interconnect_0_audio_0_avalon_audio_slave_writedata,  --                   .writedata
			readdata    => mm_interconnect_0_audio_0_avalon_audio_slave_readdata,   --                   .readdata
			irq         => open,                                                    --          interrupt.irq
			AUD_ADCDAT  => audio_0_external_interface_ADCDAT,                       -- external_interface.export
			AUD_ADCLRCK => audio_0_external_interface_ADCLRCK,                      --                   .export
			AUD_BCLK    => audio_0_external_interface_BCLK,                         --                   .export
			AUD_DACDAT  => audio_0_external_interface_DACDAT,                       --                   .export
			AUD_DACLRCK => audio_0_external_interface_DACLRCK                       --                   .export
		);

	cpu : component nios2_system_v0_cpu
		port map (
			clk                                 => clk_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,      --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,            --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                              --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	i2c_0 : component altera_avalon_i2c
		generic map (
			USE_AV_ST       => 0,
			FIFO_DEPTH      => 4,
			FIFO_DEPTH_LOG2 => 2
		)
		port map (
			clk       => clk_clk,                                      --            clock.clk
			rst_n     => rst_controller_001_reset_out_reset_ports_inv, --       reset_sink.reset_n
			intr      => open,                                         -- interrupt_sender.irq
			addr      => mm_interconnect_0_i2c_0_csr_address,          --              csr.address
			read      => mm_interconnect_0_i2c_0_csr_read,             --                 .read
			write     => mm_interconnect_0_i2c_0_csr_write,            --                 .write
			writedata => mm_interconnect_0_i2c_0_csr_writedata,        --                 .writedata
			readdata  => mm_interconnect_0_i2c_0_csr_readdata,         --                 .readdata
			sda_in    => I2C_SERIAL_SDA_IN_net,                      --       i2c_serial.sda_in
			scl_in    => I2C_SERIAL_SCL_IN_net,                      --                 .scl_in
			sda_oe    => I2C_SERIAL_SDA_OE_net,                      --                 .sda_oe
			scl_oe    => I2C_SERIAL_SCL_OE_net,                      --                 .scl_oe
			src_data  => open,                                         --      (terminated)
			src_valid => open,                                         --      (terminated)
			src_ready => '0',                                          --      (terminated)
			snk_data  => "0000000000000000",                           --      (terminated)
			snk_valid => '0',                                          --      (terminated)
			snk_ready => open                                          --      (terminated)
		);

	jtag_uart : component nios2_system_v0_jtag_uart
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	led_pio : component nios2_system_v0_led_pio
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_led_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_pio_s1_readdata,        --                    .readdata
			out_port   => led_pio_external_connection_export            -- external_connection.export
		);

	onchip_mem : component nios2_system_v0_onchip_mem
		port map (
			clk        => clk_clk,                                    --   clk1.clk
			address    => mm_interconnect_0_onchip_mem_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_mem_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_mem_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_mem_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_mem_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_mem_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_mem_s1_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,         -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req,     --       .reset_req
			freeze     => '0'                                         -- (terminated)
		);

	pll_0 : component nios2_system_v0_pll_0
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_0_outclk0_clk,       -- outclk0.clk
			locked   => open                     --  locked.export
		);

	seg_pio_0 : component nios2_system_v0_led_pio
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_seg_pio_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_seg_pio_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_seg_pio_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_seg_pio_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_seg_pio_0_s1_readdata,        --                    .readdata
			out_port   => seg_pio_0_external_connection_export            -- external_connection.export
		);

	seg_pio_1 : component nios2_system_v0_led_pio
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_seg_pio_1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_seg_pio_1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_seg_pio_1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_seg_pio_1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_seg_pio_1_s1_readdata,        --                    .readdata
			out_port   => seg_pio_1_external_connection_export            -- external_connection.export
		);

	seg_pio_2 : component nios2_system_v0_led_pio
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_seg_pio_2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_seg_pio_2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_seg_pio_2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_seg_pio_2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_seg_pio_2_s1_readdata,        --                    .readdata
			out_port   => seg_pio_2_external_connection_export            -- external_connection.export
		);

	sw_pio : component nios2_system_v0_sw_pio
		port map (
			clk      => clk_clk,                                      --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_sw_pio_s1_address,          --                  s1.address
			readdata => mm_interconnect_0_sw_pio_s1_readdata,         --                    .readdata
			in_port  => sw_pio_external_connection_export             -- external_connection.export
		);

	sys_clk_timer : component nios2_system_v0_sys_clk_timer
		port map (
			clk        => clk_clk,                                            --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,       -- reset.reset_n
			address    => mm_interconnect_0_sys_clk_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_sys_clk_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_sys_clk_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_sys_clk_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_sys_clk_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                            --   irq.irq
		);

	sysid : component nios2_system_v0_sysid
		port map (
			clock    => clk_clk,                                          --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,     --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component nios2_system_v0_mm_interconnect_0
		port map (
			clk_0_clk_clk                             => clk_clk,                                                   --                           clk_0_clk.clk
			pll_0_outclk0_clk                         => pll_0_outclk0_clk,                                         --                       pll_0_outclk0.clk
			audio_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                            -- audio_0_reset_reset_bridge_in_reset.reset
			cpu_reset_reset_bridge_in_reset_reset     => rst_controller_001_reset_out_reset,                        --     cpu_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                   => cpu_data_master_address,                                   --                     cpu_data_master.address
			cpu_data_master_waitrequest               => cpu_data_master_waitrequest,                               --                                    .waitrequest
			cpu_data_master_byteenable                => cpu_data_master_byteenable,                                --                                    .byteenable
			cpu_data_master_read                      => cpu_data_master_read,                                      --                                    .read
			cpu_data_master_readdata                  => cpu_data_master_readdata,                                  --                                    .readdata
			cpu_data_master_write                     => cpu_data_master_write,                                     --                                    .write
			cpu_data_master_writedata                 => cpu_data_master_writedata,                                 --                                    .writedata
			cpu_data_master_debugaccess               => cpu_data_master_debugaccess,                               --                                    .debugaccess
			cpu_instruction_master_address            => cpu_instruction_master_address,                            --              cpu_instruction_master.address
			cpu_instruction_master_waitrequest        => cpu_instruction_master_waitrequest,                        --                                    .waitrequest
			cpu_instruction_master_read               => cpu_instruction_master_read,                               --                                    .read
			cpu_instruction_master_readdata           => cpu_instruction_master_readdata,                           --                                    .readdata
			cpu_instruction_master_readdatavalid      => cpu_instruction_master_readdatavalid,                      --                                    .readdatavalid
			audio_0_avalon_audio_slave_address        => mm_interconnect_0_audio_0_avalon_audio_slave_address,      --          audio_0_avalon_audio_slave.address
			audio_0_avalon_audio_slave_write          => mm_interconnect_0_audio_0_avalon_audio_slave_write,        --                                    .write
			audio_0_avalon_audio_slave_read           => mm_interconnect_0_audio_0_avalon_audio_slave_read,         --                                    .read
			audio_0_avalon_audio_slave_readdata       => mm_interconnect_0_audio_0_avalon_audio_slave_readdata,     --                                    .readdata
			audio_0_avalon_audio_slave_writedata      => mm_interconnect_0_audio_0_avalon_audio_slave_writedata,    --                                    .writedata
			audio_0_avalon_audio_slave_chipselect     => mm_interconnect_0_audio_0_avalon_audio_slave_chipselect,   --                                    .chipselect
			cpu_debug_mem_slave_address               => mm_interconnect_0_cpu_debug_mem_slave_address,             --                 cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write                 => mm_interconnect_0_cpu_debug_mem_slave_write,               --                                    .write
			cpu_debug_mem_slave_read                  => mm_interconnect_0_cpu_debug_mem_slave_read,                --                                    .read
			cpu_debug_mem_slave_readdata              => mm_interconnect_0_cpu_debug_mem_slave_readdata,            --                                    .readdata
			cpu_debug_mem_slave_writedata             => mm_interconnect_0_cpu_debug_mem_slave_writedata,           --                                    .writedata
			cpu_debug_mem_slave_byteenable            => mm_interconnect_0_cpu_debug_mem_slave_byteenable,          --                                    .byteenable
			cpu_debug_mem_slave_waitrequest           => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,         --                                    .waitrequest
			cpu_debug_mem_slave_debugaccess           => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,         --                                    .debugaccess
			i2c_0_csr_address                         => mm_interconnect_0_i2c_0_csr_address,                       --                           i2c_0_csr.address
			i2c_0_csr_write                           => mm_interconnect_0_i2c_0_csr_write,                         --                                    .write
			i2c_0_csr_read                            => mm_interconnect_0_i2c_0_csr_read,                          --                                    .read
			i2c_0_csr_readdata                        => mm_interconnect_0_i2c_0_csr_readdata,                      --                                    .readdata
			i2c_0_csr_writedata                       => mm_interconnect_0_i2c_0_csr_writedata,                     --                                    .writedata
			jtag_uart_avalon_jtag_slave_address       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --         jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                    .write
			jtag_uart_avalon_jtag_slave_read          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                    .read
			jtag_uart_avalon_jtag_slave_readdata      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                    .readdata
			jtag_uart_avalon_jtag_slave_writedata     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                    .writedata
			jtag_uart_avalon_jtag_slave_waitrequest   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                    .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                    .chipselect
			led_pio_s1_address                        => mm_interconnect_0_led_pio_s1_address,                      --                          led_pio_s1.address
			led_pio_s1_write                          => mm_interconnect_0_led_pio_s1_write,                        --                                    .write
			led_pio_s1_readdata                       => mm_interconnect_0_led_pio_s1_readdata,                     --                                    .readdata
			led_pio_s1_writedata                      => mm_interconnect_0_led_pio_s1_writedata,                    --                                    .writedata
			led_pio_s1_chipselect                     => mm_interconnect_0_led_pio_s1_chipselect,                   --                                    .chipselect
			onchip_mem_s1_address                     => mm_interconnect_0_onchip_mem_s1_address,                   --                       onchip_mem_s1.address
			onchip_mem_s1_write                       => mm_interconnect_0_onchip_mem_s1_write,                     --                                    .write
			onchip_mem_s1_readdata                    => mm_interconnect_0_onchip_mem_s1_readdata,                  --                                    .readdata
			onchip_mem_s1_writedata                   => mm_interconnect_0_onchip_mem_s1_writedata,                 --                                    .writedata
			onchip_mem_s1_byteenable                  => mm_interconnect_0_onchip_mem_s1_byteenable,                --                                    .byteenable
			onchip_mem_s1_chipselect                  => mm_interconnect_0_onchip_mem_s1_chipselect,                --                                    .chipselect
			onchip_mem_s1_clken                       => mm_interconnect_0_onchip_mem_s1_clken,                     --                                    .clken
			seg_pio_0_s1_address                      => mm_interconnect_0_seg_pio_0_s1_address,                    --                        seg_pio_0_s1.address
			seg_pio_0_s1_write                        => mm_interconnect_0_seg_pio_0_s1_write,                      --                                    .write
			seg_pio_0_s1_readdata                     => mm_interconnect_0_seg_pio_0_s1_readdata,                   --                                    .readdata
			seg_pio_0_s1_writedata                    => mm_interconnect_0_seg_pio_0_s1_writedata,                  --                                    .writedata
			seg_pio_0_s1_chipselect                   => mm_interconnect_0_seg_pio_0_s1_chipselect,                 --                                    .chipselect
			seg_pio_1_s1_address                      => mm_interconnect_0_seg_pio_1_s1_address,                    --                        seg_pio_1_s1.address
			seg_pio_1_s1_write                        => mm_interconnect_0_seg_pio_1_s1_write,                      --                                    .write
			seg_pio_1_s1_readdata                     => mm_interconnect_0_seg_pio_1_s1_readdata,                   --                                    .readdata
			seg_pio_1_s1_writedata                    => mm_interconnect_0_seg_pio_1_s1_writedata,                  --                                    .writedata
			seg_pio_1_s1_chipselect                   => mm_interconnect_0_seg_pio_1_s1_chipselect,                 --                                    .chipselect
			seg_pio_2_s1_address                      => mm_interconnect_0_seg_pio_2_s1_address,                    --                        seg_pio_2_s1.address
			seg_pio_2_s1_write                        => mm_interconnect_0_seg_pio_2_s1_write,                      --                                    .write
			seg_pio_2_s1_readdata                     => mm_interconnect_0_seg_pio_2_s1_readdata,                   --                                    .readdata
			seg_pio_2_s1_writedata                    => mm_interconnect_0_seg_pio_2_s1_writedata,                  --                                    .writedata
			seg_pio_2_s1_chipselect                   => mm_interconnect_0_seg_pio_2_s1_chipselect,                 --                                    .chipselect
			sw_pio_s1_address                         => mm_interconnect_0_sw_pio_s1_address,                       --                           sw_pio_s1.address
			sw_pio_s1_readdata                        => mm_interconnect_0_sw_pio_s1_readdata,                      --                                    .readdata
			sys_clk_timer_s1_address                  => mm_interconnect_0_sys_clk_timer_s1_address,                --                    sys_clk_timer_s1.address
			sys_clk_timer_s1_write                    => mm_interconnect_0_sys_clk_timer_s1_write,                  --                                    .write
			sys_clk_timer_s1_readdata                 => mm_interconnect_0_sys_clk_timer_s1_readdata,               --                                    .readdata
			sys_clk_timer_s1_writedata                => mm_interconnect_0_sys_clk_timer_s1_writedata,              --                                    .writedata
			sys_clk_timer_s1_chipselect               => mm_interconnect_0_sys_clk_timer_s1_chipselect,             --                                    .chipselect
			sysid_control_slave_address               => mm_interconnect_0_sysid_control_slave_address,             --                 sysid_control_slave.address
			sysid_control_slave_readdata              => mm_interconnect_0_sysid_control_slave_readdata             --                                    .readdata
		);

	irq_mapper : component nios2_system_v0_irq_mapper
		port map (
			clk           => clk_clk,                            --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			sender_irq    => cpu_irq_irq                         --    sender.irq
		);

	rst_controller : component nios2_system_v0_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => pll_0_outclk0_clk,              --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component nios2_system_v0_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_sys_clk_timer_s1_write_ports_inv <= not mm_interconnect_0_sys_clk_timer_s1_write;

	mm_interconnect_0_led_pio_s1_write_ports_inv <= not mm_interconnect_0_led_pio_s1_write;

	mm_interconnect_0_seg_pio_0_s1_write_ports_inv <= not mm_interconnect_0_seg_pio_0_s1_write;

	mm_interconnect_0_seg_pio_1_s1_write_ports_inv <= not mm_interconnect_0_seg_pio_1_s1_write;

	mm_interconnect_0_seg_pio_2_s1_write_ports_inv <= not mm_interconnect_0_seg_pio_2_s1_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	audio_xclk_clk <= pll_0_outclk0_clk;
	
	I2C_SERIAL_SDA_IN_net <= i2c_0_i2c_serial_sda_inout;
	i2c_0_i2c_serial_sda_inout <= '0' when I2C_SERIAL_SDA_OE_net = '1' else 'Z';
	
	I2C_SERIAL_SCL_IN_net <= i2c_0_i2c_serial_scl_inout;
	i2c_0_i2c_serial_scl_inout <= '0' when I2C_SERIAL_SCL_OE_net = '1' else 'Z';

end architecture rtl; -- of nios2_system_v0
